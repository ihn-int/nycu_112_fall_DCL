`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Dept. of Computer Science, National Chiao Tung University
// Engineer: Chun-Jen Tsai
// 
// Create Date: 2017/05/08 15:29:41
// Design Name: 
// Module Name: lab6
// Project Name: 
// Target Devices: 
// Tool Versions:
// Description: The sample top module of lab 6: sd card reader. The behavior of
//              this module is as follows
//              1. When the SD card is initialized, display a message on the LCD.
//                 If the initialization fails, an error message will be shown.
//              2. The user can then press usr_btn[2] to trigger the sd card
//                 controller to read the super block of the sd card (located at
//                 block # 8192) into the SRAM memory.
//              3. During SD card reading time, the four LED lights will be turned on.
//                 They will be turned off when the reading is done.
//              4. The LCD will then displayer the sector just been read, and the
//                 first byte of the sector.
//              5. Everytime you press usr_btn[2], the next byte will be displayed.
// 
// Dependencies: clk_divider, LCD_module, debounce, sd_card
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module lab8(
  // General system I/O ports
  input  clk,
  input  reset_n,
  input  [3:0] usr_btn,
  output [3:0] usr_led,

  // SD card specific I/O ports
  output spi_ss,
  output spi_sck,
  output spi_mosi,
  input  spi_miso,

  // 1602 LCD Module Interface
  output LCD_RS,
  output LCD_RW,
  output LCD_E,
  output [3:0] LCD_D
);

localparam [2:0] S_MAIN_INIT = 3'b000, S_MAIN_IDLE = 3'b001,
                 S_MAIN_WAIT = 3'b010, S_MAIN_FIND = 3'b011,
                 S_MAIN_READ = 3'b100, S_MAIN_NBLK = 3'b101,
                 S_MAIN_DONE = 3'b110;

// Declare system variables
wire btn_level, btn_pressed;
reg  prev_btn_level;
reg  [2:0] P, P_next;
reg  [9:0] sd_counter;

reg  [127:0] row_A = "SD card cannot  ";
reg  [127:0] row_B = "be initialized! ";
reg  done_flag; // Signals the completion of reading one SD sector.

// Declare SD card interface signals
wire clk_sel;
wire clk_500k;
reg  rd_req;
reg  [31:0] rd_addr;
wire init_finished;
wire [7:0] sd_dout;
wire sd_valid;

assign clk_sel = (init_finished)? clk : clk_500k; // clock for the SD controller
assign usr_led = P;

reg[63:0] volc;
reg[15:0] cnt;
reg[2:0] word_cnt;


clk_divider#(200) clk_divider0(
  .clk(clk),
  .reset(~reset_n),
  .clk_out(clk_500k)
);

debounce btn_db0(
  .clk(clk),
  .btn_input(usr_btn[2]),
  .btn_output(btn_level)
);

LCD_module lcd0( 
  .clk(clk),
  .reset(~reset_n),
  .row_A(row_A),
  .row_B(row_B),
  .LCD_E(LCD_E),
  .LCD_RS(LCD_RS),
  .LCD_RW(LCD_RW),
  .LCD_D(LCD_D)
);

sd_card sd_card0(
  .cs(spi_ss),
  .sclk(spi_sck),
  .mosi(spi_mosi),
  .miso(spi_miso),

  .clk(clk_sel),
  .rst(~reset_n),
  .rd_req(rd_req),
  .block_addr(rd_addr),
  .init_finished(init_finished),
  .dout(sd_dout),
  .sd_valid(sd_valid)
);

//
// Enable one cycle of btn_pressed per each button hit
//
always @(posedge clk) begin
  if (~reset_n)
    prev_btn_level <= 0;
  else
    prev_btn_level <= btn_level;
end

assign btn_pressed = (btn_level == 1 && prev_btn_level == 0)? 1 : 0;

// ------------------------------------------------------------------------
// FSM of the SD card reader that reads the super block (512 bytes)
always @(posedge clk) begin
  if (~reset_n) begin
    P <= S_MAIN_INIT;
  end
  else begin
    P <= P_next;
  end
end

always @(*) begin // FSM next-state logic
  case (P)
    S_MAIN_INIT: // wait for SD card initialization
      if (init_finished == 1) P_next = S_MAIN_IDLE;
      else P_next = S_MAIN_INIT;
    S_MAIN_IDLE: // wait for button click
      if (btn_pressed == 1) P_next = S_MAIN_WAIT;
      else P_next = S_MAIN_IDLE;
    S_MAIN_WAIT: // issue a rd_req to the SD controller until it's ready
      P_next = S_MAIN_FIND;
    S_MAIN_FIND: // find the tag
      if(volc == "DLAB_TAG") P_next = S_MAIN_READ;
      else if(sd_counter == 512) P_next = S_MAIN_WAIT;
      else P_next = S_MAIN_FIND;
    S_MAIN_READ: // wait for the input data to enter the SRAM buffer
      if (sd_counter == 512) P_next = S_MAIN_NBLK;
      else if (volc == "DLAB_END") P_next = S_MAIN_DONE;
      else P_next = S_MAIN_READ;
    S_MAIN_NBLK: //
      P_next = S_MAIN_READ;
    S_MAIN_DONE: // read byte 0 of the superblock from sram[]
      P_next = S_MAIN_DONE;
    default:
      P_next = S_MAIN_IDLE;
  endcase
end

// FSM output logic: controls the 'rd_req' and 'rd_addr' signals.
always @(*) begin
  rd_req = (P == S_MAIN_WAIT) || (P == S_MAIN_NBLK);
  
end

always @(posedge clk) begin
  if (~reset_n) rd_addr <= 32'h2000;
  else if ((P == S_MAIN_WAIT) || (P == S_MAIN_NBLK)) rd_addr <= rd_addr + 1;
   // In lab 6, change this line to scan all blocks
end

// FSM output logic: controls the 'sd_counter' signal.
// SD card read address incrementer
always @(posedge clk) begin
  if (~reset_n || P == S_MAIN_WAIT || P == S_MAIN_NBLK)
    sd_counter <= 0;
  else if ((P == S_MAIN_FIND  || P == S_MAIN_READ ) && sd_valid)
    sd_counter <= sd_counter + 1;
end

always@(posedge clk) begin
  if(~reset_n) volc = 64'h0;
  else if(sd_valid && (P == S_MAIN_FIND || P == S_MAIN_READ)) begin
    volc <= { volc[55:0] , sd_dout};
  end
end

always@(posedge clk) begin
  if(~reset_n) begin
    cnt = 0;
    word_cnt = 0;
  end
  else if(P == S_MAIN_READ && sd_valid) begin
    if((sd_dout >= "A" && sd_dout <= "Z") ||
       (sd_dout >= "a" && sd_dout <= "z"))
      word_cnt <= (word_cnt[2]) ? 4 : word_cnt + 1;
    else begin
      if(word_cnt == 3) cnt <= cnt + 1;
      word_cnt <= 0;    
    end
  end
end

// End of the FSM of the SD card reader
// ------------------------------------------------------------------------

// ------------------------------------------------------------------------
// LCD Display function.
always @(posedge clk) begin
  if (~reset_n) begin
    row_A = "SD card cannot  ";
    row_B = "be initialized! ";
  end else if (P == S_MAIN_DONE) begin
    row_A <= { "Found ",
               ((cnt[15:12] > 9) ? "7" : "0") + cnt[15:12],
               ((cnt[11: 8] > 9) ? "7" : "0") + cnt[11: 8],
               ((cnt[7 : 4] > 9) ? "7" : "0") + cnt[7 : 4],
               ((cnt[3 : 0] > 9) ? "7" : "0") + cnt[3 : 0],
               " words"
             };
    row_B <= "in the text file";
  end
  else if (P == S_MAIN_IDLE) begin
    row_A <= "Hit BTN2 to read";
    row_B <= "the SD card ... ";
  end
end
// End of the LCD display function
// ------------------------------------------------------------------------

endmodule
